ENTITY aula_3 IS
    PORT (
        SW : IN bit_vector(9 DOWNTO 0);
        HEX0 : OUT bit_vector(6 DOWNTO 0);
        HEX1 : OUT bit_vector(6 DOWNTO 0);
        HEX2 : OUT bit_vector(6 DOWNTO 0);
        HEX3 : OUT bit_vector(6 DOWNTO 0);
        HEX4 : OUT bit_vector(6 DOWNTO 0);
        HEX5 : OUT bit_vector(6 DOWNTO 0)
    );
END aula_3;